magic
tech sky130A
magscale 1 2
timestamp 1729221706
<< nmos >>
rect -286 109 -86 509
rect 86 109 286 509
rect -286 -509 -86 -109
rect 86 -509 286 -109
<< ndiff >>
rect -344 497 -286 509
rect -344 121 -332 497
rect -298 121 -286 497
rect -344 109 -286 121
rect -86 497 -28 509
rect -86 121 -74 497
rect -40 121 -28 497
rect -86 109 -28 121
rect 28 497 86 509
rect 28 121 40 497
rect 74 121 86 497
rect 28 109 86 121
rect 286 497 344 509
rect 286 121 298 497
rect 332 121 344 497
rect 286 109 344 121
rect -344 -121 -286 -109
rect -344 -497 -332 -121
rect -298 -497 -286 -121
rect -344 -509 -286 -497
rect -86 -121 -28 -109
rect -86 -497 -74 -121
rect -40 -497 -28 -121
rect -86 -509 -28 -497
rect 28 -121 86 -109
rect 28 -497 40 -121
rect 74 -497 86 -121
rect 28 -509 86 -497
rect 286 -121 344 -109
rect 286 -497 298 -121
rect 332 -497 344 -121
rect 286 -509 344 -497
<< ndiffc >>
rect -332 121 -298 497
rect -74 121 -40 497
rect 40 121 74 497
rect 298 121 332 497
rect -332 -497 -298 -121
rect -74 -497 -40 -121
rect 40 -497 74 -121
rect 298 -497 332 -121
<< poly >>
rect -286 581 -86 597
rect -286 547 -270 581
rect -102 547 -86 581
rect -286 509 -86 547
rect 86 581 286 597
rect 86 547 102 581
rect 270 547 286 581
rect 86 509 286 547
rect -286 71 -86 109
rect -286 37 -270 71
rect -102 37 -86 71
rect -286 21 -86 37
rect 86 71 286 109
rect 86 37 102 71
rect 270 37 286 71
rect 86 21 286 37
rect -286 -37 -86 -21
rect -286 -71 -270 -37
rect -102 -71 -86 -37
rect -286 -109 -86 -71
rect 86 -37 286 -21
rect 86 -71 102 -37
rect 270 -71 286 -37
rect 86 -109 286 -71
rect -286 -547 -86 -509
rect -286 -581 -270 -547
rect -102 -581 -86 -547
rect -286 -597 -86 -581
rect 86 -547 286 -509
rect 86 -581 102 -547
rect 270 -581 286 -547
rect 86 -597 286 -581
<< polycont >>
rect -270 547 -102 581
rect 102 547 270 581
rect -270 37 -102 71
rect 102 37 270 71
rect -270 -71 -102 -37
rect 102 -71 270 -37
rect -270 -581 -102 -547
rect 102 -581 270 -547
<< locali >>
rect -286 547 -270 581
rect -102 547 -86 581
rect 86 547 102 581
rect 270 547 286 581
rect -332 497 -298 513
rect -332 105 -298 121
rect -74 497 -40 513
rect -74 105 -40 121
rect 40 497 74 513
rect 40 105 74 121
rect 298 497 332 513
rect 298 105 332 121
rect -286 37 -270 71
rect -102 37 -86 71
rect 86 37 102 71
rect 270 37 286 71
rect -286 -71 -270 -37
rect -102 -71 -86 -37
rect 86 -71 102 -37
rect 270 -71 286 -37
rect -332 -121 -298 -105
rect -332 -513 -298 -497
rect -74 -121 -40 -105
rect -74 -513 -40 -497
rect 40 -121 74 -105
rect 40 -513 74 -497
rect 298 -121 332 -105
rect 298 -513 332 -497
rect -286 -581 -270 -547
rect -102 -581 -86 -547
rect 86 -581 102 -547
rect 270 -581 286 -547
<< viali >>
rect -249 547 -123 581
rect 123 547 249 581
rect -332 121 -298 497
rect -74 121 -40 497
rect 40 121 74 497
rect 298 121 332 497
rect -249 37 -123 71
rect 123 37 249 71
rect -249 -71 -123 -37
rect 123 -71 249 -37
rect -332 -497 -298 -121
rect -74 -497 -40 -121
rect 40 -497 74 -121
rect 298 -497 332 -121
rect -249 -581 -123 -547
rect 123 -581 249 -547
<< metal1 >>
rect -261 581 -111 587
rect -261 547 -249 581
rect -123 547 -111 581
rect -261 541 -111 547
rect 111 581 261 587
rect 111 547 123 581
rect 249 547 261 581
rect 111 541 261 547
rect -338 497 -292 509
rect -338 121 -332 497
rect -298 121 -292 497
rect -338 109 -292 121
rect -80 497 -34 509
rect -80 121 -74 497
rect -40 121 -34 497
rect -80 109 -34 121
rect 34 497 80 509
rect 34 121 40 497
rect 74 121 80 497
rect 34 109 80 121
rect 292 497 338 509
rect 292 121 298 497
rect 332 121 338 497
rect 292 109 338 121
rect -261 71 -111 77
rect -261 37 -249 71
rect -123 37 -111 71
rect -261 31 -111 37
rect 111 71 261 77
rect 111 37 123 71
rect 249 37 261 71
rect 111 31 261 37
rect -261 -37 -111 -31
rect -261 -71 -249 -37
rect -123 -71 -111 -37
rect -261 -77 -111 -71
rect 111 -37 261 -31
rect 111 -71 123 -37
rect 249 -71 261 -37
rect 111 -77 261 -71
rect -338 -121 -292 -109
rect -338 -497 -332 -121
rect -298 -497 -292 -121
rect -338 -509 -292 -497
rect -80 -121 -34 -109
rect -80 -497 -74 -121
rect -40 -497 -34 -121
rect -80 -509 -34 -497
rect 34 -121 80 -109
rect 34 -497 40 -121
rect 74 -497 80 -121
rect 34 -509 80 -497
rect 292 -121 338 -109
rect 292 -497 298 -121
rect 332 -497 338 -121
rect 292 -509 338 -497
rect -261 -547 -111 -541
rect -261 -581 -249 -547
rect -123 -581 -111 -547
rect -261 -587 -111 -581
rect 111 -547 261 -541
rect 111 -581 123 -547
rect 249 -581 261 -547
rect 111 -587 261 -581
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 1 m 2 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 0 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
