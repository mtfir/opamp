magic
tech sky130A
magscale 1 2
timestamp 1729406401
<< nwell >>
rect -228 -89 874 2597
<< nsubdiff >>
rect -192 2527 -132 2561
rect 778 2527 838 2561
rect -192 2501 -158 2527
rect 804 2501 838 2527
rect -192 -19 -158 7
rect 804 -19 838 7
rect -192 -53 -132 -19
rect 778 -53 838 -19
<< nsubdiffcont >>
rect -132 2527 778 2561
rect -192 7 -158 2501
rect 804 7 838 2501
rect -132 -53 778 -19
<< poly >>
rect 94 640 294 2505
rect 352 3 552 1869
<< locali >>
rect -192 2527 -132 2561
rect 778 2527 838 2561
rect -192 2501 -158 2527
rect -192 -19 -158 7
rect 804 2501 838 2527
rect 804 -19 838 7
rect -192 -53 -132 -19
rect 778 -53 838 -19
<< viali >>
rect 626 2527 676 2561
rect -30 -53 20 -19
<< metal1 >>
rect 614 2561 688 2567
rect 614 2527 626 2561
rect 676 2527 688 2561
rect -42 2408 32 2495
rect 377 2408 527 2495
rect 614 2408 688 2527
rect -98 2384 88 2408
rect -111 2008 -101 2384
rect -49 2008 88 2384
rect 300 2008 744 2408
rect -42 1772 32 1859
rect -98 1760 88 1772
rect -98 1384 39 1760
rect 91 1384 101 1760
rect -98 1372 88 1384
rect -98 1124 88 1136
rect -98 748 39 1124
rect 91 748 101 1124
rect -98 736 88 748
rect -42 695 32 736
rect -42 649 269 695
rect 300 500 346 2008
rect 377 1813 688 1859
rect 614 1772 688 1813
rect 558 1760 744 1772
rect 545 1384 555 1760
rect 607 1384 744 1760
rect 558 1372 744 1384
rect 558 1124 744 1136
rect 545 748 555 1124
rect 607 748 744 1124
rect 558 736 744 748
rect 614 649 688 736
rect -98 100 346 500
rect 558 488 744 500
rect 558 112 695 488
rect 747 112 757 488
rect 558 100 744 112
rect -42 -19 32 100
rect 119 14 269 100
rect 614 13 688 100
rect -42 -53 -30 -19
rect 20 -53 32 -19
rect -42 -59 32 -53
<< via1 >>
rect -101 2008 -49 2384
rect 39 1384 91 1760
rect 39 748 91 1124
rect 555 1384 607 1760
rect 555 748 607 1124
rect 695 112 747 488
<< metal2 >>
rect -101 2384 -49 2394
rect -101 1916 -49 2008
rect -101 1864 747 1916
rect -101 644 -49 1864
rect 39 1760 91 1770
rect 39 1280 91 1384
rect 553 1760 609 1770
rect 553 1374 609 1384
rect 39 1228 607 1280
rect 37 1124 93 1134
rect 37 738 93 748
rect 555 1124 607 1228
rect 555 738 607 748
rect 695 644 747 1864
rect -101 592 747 644
rect 695 488 747 592
rect 695 102 747 112
<< via2 >>
rect 553 1384 555 1760
rect 555 1384 607 1760
rect 607 1384 609 1760
rect 37 748 39 1124
rect 39 748 91 1124
rect 91 748 93 1124
<< metal3 >>
rect 543 1760 619 1765
rect 543 1384 553 1760
rect 609 1384 619 1760
rect 543 1292 619 1384
rect 27 1216 619 1292
rect 27 1124 103 1216
rect 27 748 37 1124
rect 93 748 103 1124
rect 27 743 103 748
use sky130_fd_pr__pfet_01v8_EZH3Y7  sky130_fd_pr__pfet_01v8_EZH3Y7_0
timestamp 1729184099
transform 1 0 651 0 1 1254
box -135 -1254 135 1254
use sky130_fd_pr__pfet_01v8_EZH3Y7  sky130_fd_pr__pfet_01v8_EZH3Y7_1
timestamp 1729184099
transform 1 0 -5 0 1 1254
box -135 -1254 135 1254
use sky130_fd_pr__pfet_01v8_SD2LB7  sky130_fd_pr__pfet_01v8_SD2LB7_0
timestamp 1729184099
transform 1 0 323 0 1 1254
box -323 -1254 323 1254
<< labels >>
flabel metal1 448 2223 449 2224 0 FreeSans 160 0 0 0 VDD
port 0 nsew
flabel metal1 -10 2214 -9 2215 0 FreeSans 160 0 0 0 D5
port 1 nsew
flabel metal1 -8 1587 -8 1587 0 FreeSans 160 0 0 0 D1
port 2 nsew
flabel metal1 -12 960 -12 960 0 FreeSans 160 0 0 0 D2
port 3 nsew
<< end >>
