magic
tech sky130A
magscale 1 2
timestamp 1729184099
<< error_p >>
rect -135 654 135 872
rect -135 18 135 236
rect -135 -618 135 -400
<< nwell >>
rect -135 654 135 1254
rect -135 18 135 618
rect -135 -618 135 -18
rect -135 -1254 135 -654
<< pmos >>
rect -41 754 41 1154
rect -41 118 41 518
rect -41 -518 41 -118
rect -41 -1154 41 -754
<< pdiff >>
rect -99 1142 -41 1154
rect -99 766 -87 1142
rect -53 766 -41 1142
rect -99 754 -41 766
rect 41 1142 99 1154
rect 41 766 53 1142
rect 87 766 99 1142
rect 41 754 99 766
rect -99 506 -41 518
rect -99 130 -87 506
rect -53 130 -41 506
rect -99 118 -41 130
rect 41 506 99 518
rect 41 130 53 506
rect 87 130 99 506
rect 41 118 99 130
rect -99 -130 -41 -118
rect -99 -506 -87 -130
rect -53 -506 -41 -130
rect -99 -518 -41 -506
rect 41 -130 99 -118
rect 41 -506 53 -130
rect 87 -506 99 -130
rect 41 -518 99 -506
rect -99 -766 -41 -754
rect -99 -1142 -87 -766
rect -53 -1142 -41 -766
rect -99 -1154 -41 -1142
rect 41 -766 99 -754
rect 41 -1142 53 -766
rect 87 -1142 99 -766
rect 41 -1154 99 -1142
<< pdiffc >>
rect -87 766 -53 1142
rect 53 766 87 1142
rect -87 130 -53 506
rect 53 130 87 506
rect -87 -506 -53 -130
rect 53 -506 87 -130
rect -87 -1142 -53 -766
rect 53 -1142 87 -766
<< poly >>
rect -41 1235 41 1251
rect -41 1201 -25 1235
rect 25 1201 41 1235
rect -41 1154 41 1201
rect -41 707 41 754
rect -41 673 -25 707
rect 25 673 41 707
rect -41 657 41 673
rect -41 599 41 615
rect -41 565 -25 599
rect 25 565 41 599
rect -41 518 41 565
rect -41 71 41 118
rect -41 37 -25 71
rect 25 37 41 71
rect -41 21 41 37
rect -41 -37 41 -21
rect -41 -71 -25 -37
rect 25 -71 41 -37
rect -41 -118 41 -71
rect -41 -565 41 -518
rect -41 -599 -25 -565
rect 25 -599 41 -565
rect -41 -615 41 -599
rect -41 -673 41 -657
rect -41 -707 -25 -673
rect 25 -707 41 -673
rect -41 -754 41 -707
rect -41 -1201 41 -1154
rect -41 -1235 -25 -1201
rect 25 -1235 41 -1201
rect -41 -1251 41 -1235
<< polycont >>
rect -25 1201 25 1235
rect -25 673 25 707
rect -25 565 25 599
rect -25 37 25 71
rect -25 -71 25 -37
rect -25 -599 25 -565
rect -25 -707 25 -673
rect -25 -1235 25 -1201
<< locali >>
rect -41 1201 -25 1235
rect 25 1201 41 1235
rect -87 1142 -53 1158
rect -87 750 -53 766
rect 53 1142 87 1158
rect 53 750 87 766
rect -41 673 -25 707
rect 25 673 41 707
rect -41 565 -25 599
rect 25 565 41 599
rect -87 506 -53 522
rect -87 114 -53 130
rect 53 506 87 522
rect 53 114 87 130
rect -41 37 -25 71
rect 25 37 41 71
rect -41 -71 -25 -37
rect 25 -71 41 -37
rect -87 -130 -53 -114
rect -87 -522 -53 -506
rect 53 -130 87 -114
rect 53 -522 87 -506
rect -41 -599 -25 -565
rect 25 -599 41 -565
rect -41 -707 -25 -673
rect 25 -707 41 -673
rect -87 -766 -53 -750
rect -87 -1158 -53 -1142
rect 53 -766 87 -750
rect 53 -1158 87 -1142
rect -41 -1235 -25 -1201
rect 25 -1235 41 -1201
<< viali >>
rect -25 1201 25 1235
rect -87 766 -53 1142
rect 53 766 87 1142
rect -25 673 25 707
rect -25 565 25 599
rect -87 130 -53 506
rect 53 130 87 506
rect -25 37 25 71
rect -25 -71 25 -37
rect -87 -506 -53 -130
rect 53 -506 87 -130
rect -25 -599 25 -565
rect -25 -707 25 -673
rect -87 -1142 -53 -766
rect 53 -1142 87 -766
rect -25 -1235 25 -1201
<< metal1 >>
rect -37 1235 37 1241
rect -37 1201 -25 1235
rect 25 1201 37 1235
rect -37 1195 37 1201
rect -93 1142 -47 1154
rect -93 766 -87 1142
rect -53 766 -47 1142
rect -93 754 -47 766
rect 47 1142 93 1154
rect 47 766 53 1142
rect 87 766 93 1142
rect 47 754 93 766
rect -37 707 37 713
rect -37 673 -25 707
rect 25 673 37 707
rect -37 667 37 673
rect -37 599 37 605
rect -37 565 -25 599
rect 25 565 37 599
rect -37 559 37 565
rect -93 506 -47 518
rect -93 130 -87 506
rect -53 130 -47 506
rect -93 118 -47 130
rect 47 506 93 518
rect 47 130 53 506
rect 87 130 93 506
rect 47 118 93 130
rect -37 71 37 77
rect -37 37 -25 71
rect 25 37 37 71
rect -37 31 37 37
rect -37 -37 37 -31
rect -37 -71 -25 -37
rect 25 -71 37 -37
rect -37 -77 37 -71
rect -93 -130 -47 -118
rect -93 -506 -87 -130
rect -53 -506 -47 -130
rect -93 -518 -47 -506
rect 47 -130 93 -118
rect 47 -506 53 -130
rect 87 -506 93 -130
rect 47 -518 93 -506
rect -37 -565 37 -559
rect -37 -599 -25 -565
rect 25 -599 37 -565
rect -37 -605 37 -599
rect -37 -673 37 -667
rect -37 -707 -25 -673
rect 25 -707 37 -673
rect -37 -713 37 -707
rect -93 -766 -47 -754
rect -93 -1142 -87 -766
rect -53 -1142 -47 -766
rect -93 -1154 -47 -1142
rect 47 -766 93 -754
rect 47 -1142 53 -766
rect 87 -1142 93 -766
rect 47 -1154 93 -1142
rect -37 -1201 37 -1195
rect -37 -1235 -25 -1201
rect 25 -1235 37 -1201
rect -37 -1241 37 -1235
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 0.41 m 4 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
