magic
tech sky130A
magscale 1 2
timestamp 1729325631
<< nmos >>
rect -189 527 -29 727
rect 29 527 189 727
rect -189 109 -29 309
rect 29 109 189 309
rect -189 -309 -29 -109
rect 29 -309 189 -109
rect -189 -727 -29 -527
rect 29 -727 189 -527
<< ndiff >>
rect -247 715 -189 727
rect -247 539 -235 715
rect -201 539 -189 715
rect -247 527 -189 539
rect -29 715 29 727
rect -29 539 -17 715
rect 17 539 29 715
rect -29 527 29 539
rect 189 715 247 727
rect 189 539 201 715
rect 235 539 247 715
rect 189 527 247 539
rect -247 297 -189 309
rect -247 121 -235 297
rect -201 121 -189 297
rect -247 109 -189 121
rect -29 297 29 309
rect -29 121 -17 297
rect 17 121 29 297
rect -29 109 29 121
rect 189 297 247 309
rect 189 121 201 297
rect 235 121 247 297
rect 189 109 247 121
rect -247 -121 -189 -109
rect -247 -297 -235 -121
rect -201 -297 -189 -121
rect -247 -309 -189 -297
rect -29 -121 29 -109
rect -29 -297 -17 -121
rect 17 -297 29 -121
rect -29 -309 29 -297
rect 189 -121 247 -109
rect 189 -297 201 -121
rect 235 -297 247 -121
rect 189 -309 247 -297
rect -247 -539 -189 -527
rect -247 -715 -235 -539
rect -201 -715 -189 -539
rect -247 -727 -189 -715
rect -29 -539 29 -527
rect -29 -715 -17 -539
rect 17 -715 29 -539
rect -29 -727 29 -715
rect 189 -539 247 -527
rect 189 -715 201 -539
rect 235 -715 247 -539
rect 189 -727 247 -715
<< ndiffc >>
rect -235 539 -201 715
rect -17 539 17 715
rect 201 539 235 715
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect -235 -715 -201 -539
rect -17 -715 17 -539
rect 201 -715 235 -539
<< poly >>
rect -189 799 -29 815
rect -189 765 -173 799
rect -45 765 -29 799
rect -189 727 -29 765
rect 29 799 189 815
rect 29 765 45 799
rect 173 765 189 799
rect 29 727 189 765
rect -189 489 -29 527
rect -189 455 -173 489
rect -45 455 -29 489
rect -189 439 -29 455
rect 29 489 189 527
rect 29 455 45 489
rect 173 455 189 489
rect 29 439 189 455
rect -189 381 -29 397
rect -189 347 -173 381
rect -45 347 -29 381
rect -189 309 -29 347
rect 29 381 189 397
rect 29 347 45 381
rect 173 347 189 381
rect 29 309 189 347
rect -189 71 -29 109
rect -189 37 -173 71
rect -45 37 -29 71
rect -189 21 -29 37
rect 29 71 189 109
rect 29 37 45 71
rect 173 37 189 71
rect 29 21 189 37
rect -189 -37 -29 -21
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect -189 -109 -29 -71
rect 29 -37 189 -21
rect 29 -71 45 -37
rect 173 -71 189 -37
rect 29 -109 189 -71
rect -189 -347 -29 -309
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect -189 -397 -29 -381
rect 29 -347 189 -309
rect 29 -381 45 -347
rect 173 -381 189 -347
rect 29 -397 189 -381
rect -189 -455 -29 -439
rect -189 -489 -173 -455
rect -45 -489 -29 -455
rect -189 -527 -29 -489
rect 29 -455 189 -439
rect 29 -489 45 -455
rect 173 -489 189 -455
rect 29 -527 189 -489
rect -189 -765 -29 -727
rect -189 -799 -173 -765
rect -45 -799 -29 -765
rect -189 -815 -29 -799
rect 29 -765 189 -727
rect 29 -799 45 -765
rect 173 -799 189 -765
rect 29 -815 189 -799
<< polycont >>
rect -173 765 -45 799
rect 45 765 173 799
rect -173 455 -45 489
rect 45 455 173 489
rect -173 347 -45 381
rect 45 347 173 381
rect -173 37 -45 71
rect 45 37 173 71
rect -173 -71 -45 -37
rect 45 -71 173 -37
rect -173 -381 -45 -347
rect 45 -381 173 -347
rect -173 -489 -45 -455
rect 45 -489 173 -455
rect -173 -799 -45 -765
rect 45 -799 173 -765
<< locali >>
rect -189 765 -173 799
rect -45 765 -29 799
rect 29 765 45 799
rect 173 765 189 799
rect -235 715 -201 731
rect -235 523 -201 539
rect -17 715 17 731
rect -17 523 17 539
rect 201 715 235 731
rect 201 523 235 539
rect -189 455 -173 489
rect -45 455 -29 489
rect 29 455 45 489
rect 173 455 189 489
rect -189 347 -173 381
rect -45 347 -29 381
rect 29 347 45 381
rect 173 347 189 381
rect -235 297 -201 313
rect -235 105 -201 121
rect -17 297 17 313
rect -17 105 17 121
rect 201 297 235 313
rect 201 105 235 121
rect -189 37 -173 71
rect -45 37 -29 71
rect 29 37 45 71
rect 173 37 189 71
rect -189 -71 -173 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 173 -71 189 -37
rect -235 -121 -201 -105
rect -235 -313 -201 -297
rect -17 -121 17 -105
rect -17 -313 17 -297
rect 201 -121 235 -105
rect 201 -313 235 -297
rect -189 -381 -173 -347
rect -45 -381 -29 -347
rect 29 -381 45 -347
rect 173 -381 189 -347
rect -189 -489 -173 -455
rect -45 -489 -29 -455
rect 29 -489 45 -455
rect 173 -489 189 -455
rect -235 -539 -201 -523
rect -235 -731 -201 -715
rect -17 -539 17 -523
rect -17 -731 17 -715
rect 201 -539 235 -523
rect 201 -731 235 -715
rect -189 -799 -173 -765
rect -45 -799 -29 -765
rect 29 -799 45 -765
rect 173 -799 189 -765
<< viali >>
rect -154 765 -64 799
rect 64 765 154 799
rect -235 539 -201 715
rect -17 539 17 715
rect 201 539 235 715
rect -154 455 -64 489
rect 64 455 154 489
rect -154 347 -64 381
rect 64 347 154 381
rect -235 121 -201 297
rect -17 121 17 297
rect 201 121 235 297
rect -154 37 -64 71
rect 64 37 154 71
rect -154 -71 -64 -37
rect 64 -71 154 -37
rect -235 -297 -201 -121
rect -17 -297 17 -121
rect 201 -297 235 -121
rect -154 -381 -64 -347
rect 64 -381 154 -347
rect -154 -489 -64 -455
rect 64 -489 154 -455
rect -235 -715 -201 -539
rect -17 -715 17 -539
rect 201 -715 235 -539
rect -154 -799 -64 -765
rect 64 -799 154 -765
<< metal1 >>
rect -166 799 -52 805
rect -166 765 -154 799
rect -64 765 -52 799
rect -166 759 -52 765
rect 52 799 166 805
rect 52 765 64 799
rect 154 765 166 799
rect 52 759 166 765
rect -241 715 -195 727
rect -241 539 -235 715
rect -201 539 -195 715
rect -241 527 -195 539
rect -23 715 23 727
rect -23 539 -17 715
rect 17 539 23 715
rect -23 527 23 539
rect 195 715 241 727
rect 195 539 201 715
rect 235 539 241 715
rect 195 527 241 539
rect -166 489 -52 495
rect -166 455 -154 489
rect -64 455 -52 489
rect -166 449 -52 455
rect 52 489 166 495
rect 52 455 64 489
rect 154 455 166 489
rect 52 449 166 455
rect -166 381 -52 387
rect -166 347 -154 381
rect -64 347 -52 381
rect -166 341 -52 347
rect 52 381 166 387
rect 52 347 64 381
rect 154 347 166 381
rect 52 341 166 347
rect -241 297 -195 309
rect -241 121 -235 297
rect -201 121 -195 297
rect -241 109 -195 121
rect -23 297 23 309
rect -23 121 -17 297
rect 17 121 23 297
rect -23 109 23 121
rect 195 297 241 309
rect 195 121 201 297
rect 235 121 241 297
rect 195 109 241 121
rect -166 71 -52 77
rect -166 37 -154 71
rect -64 37 -52 71
rect -166 31 -52 37
rect 52 71 166 77
rect 52 37 64 71
rect 154 37 166 71
rect 52 31 166 37
rect -166 -37 -52 -31
rect -166 -71 -154 -37
rect -64 -71 -52 -37
rect -166 -77 -52 -71
rect 52 -37 166 -31
rect 52 -71 64 -37
rect 154 -71 166 -37
rect 52 -77 166 -71
rect -241 -121 -195 -109
rect -241 -297 -235 -121
rect -201 -297 -195 -121
rect -241 -309 -195 -297
rect -23 -121 23 -109
rect -23 -297 -17 -121
rect 17 -297 23 -121
rect -23 -309 23 -297
rect 195 -121 241 -109
rect 195 -297 201 -121
rect 235 -297 241 -121
rect 195 -309 241 -297
rect -166 -347 -52 -341
rect -166 -381 -154 -347
rect -64 -381 -52 -347
rect -166 -387 -52 -381
rect 52 -347 166 -341
rect 52 -381 64 -347
rect 154 -381 166 -347
rect 52 -387 166 -381
rect -166 -455 -52 -449
rect -166 -489 -154 -455
rect -64 -489 -52 -455
rect -166 -495 -52 -489
rect 52 -455 166 -449
rect 52 -489 64 -455
rect 154 -489 166 -455
rect 52 -495 166 -489
rect -241 -539 -195 -527
rect -241 -715 -235 -539
rect -201 -715 -195 -539
rect -241 -727 -195 -715
rect -23 -539 23 -527
rect -23 -715 -17 -539
rect 17 -715 23 -539
rect -23 -727 23 -715
rect 195 -539 241 -527
rect 195 -715 201 -539
rect 235 -715 241 -539
rect 195 -727 241 -715
rect -166 -765 -52 -759
rect -166 -799 -154 -765
rect -64 -799 -52 -765
rect -166 -805 -52 -799
rect 52 -765 166 -759
rect 52 -799 64 -765
rect 154 -799 166 -765
rect 52 -805 166 -799
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1 l 0.8 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 70 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
