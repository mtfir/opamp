magic
tech sky130A
magscale 1 2
timestamp 1729352936
<< psubdiff >>
rect -246 1661 -186 1695
rect 680 1661 740 1695
rect -246 1635 -212 1661
rect 706 1635 740 1661
rect -246 -31 -212 -5
rect 706 -31 740 -5
rect -246 -65 -186 -31
rect 680 -65 740 -31
<< psubdiffcont >>
rect -186 1661 680 1695
rect -246 -5 -212 1635
rect 706 -5 740 1635
rect -186 -65 680 -31
<< poly >>
rect 58 -1 218 1630
rect 276 0 436 1631
<< locali >>
rect -246 1661 -186 1695
rect 680 1661 740 1695
rect -246 1635 -212 1661
rect -246 -31 -212 -5
rect 706 1635 740 1661
rect 706 -31 740 -5
rect -246 -65 -186 -31
rect 680 -65 740 -31
<< viali >>
rect 230 1661 264 1695
rect 230 -65 264 -31
<< metal1 >>
rect 218 1695 276 1701
rect 218 1661 230 1695
rect 264 1661 276 1695
rect 218 1655 276 1661
rect 83 1620 93 1623
rect -96 1574 93 1620
rect -96 1542 -4 1574
rect 83 1571 93 1574
rect 183 1620 193 1623
rect 183 1574 195 1620
rect 183 1571 193 1574
rect -152 1342 52 1542
rect -96 1264 -4 1342
rect -94 1202 -84 1205
rect -96 1153 -84 1202
rect -16 1202 -6 1205
rect -16 1153 -4 1202
rect -96 1124 -4 1153
rect -152 924 52 1124
rect -96 706 -4 924
rect -152 506 52 706
rect -96 477 -4 506
rect -96 429 -84 477
rect -94 425 -84 429
rect -16 429 -4 477
rect -16 425 -6 429
rect -96 288 -4 366
rect -152 88 52 288
rect -96 56 -4 88
rect 83 56 93 59
rect -96 10 93 56
rect 83 7 93 10
rect 183 56 193 59
rect 183 10 195 56
rect 183 7 193 10
rect 224 -25 270 1655
rect 301 1571 311 1623
rect 401 1571 411 1623
rect 498 1542 590 1620
rect 442 1342 646 1542
rect 498 1313 590 1342
rect 498 1264 510 1313
rect 500 1261 510 1264
rect 578 1264 590 1313
rect 578 1261 588 1264
rect 299 1156 590 1202
rect 498 1124 590 1156
rect 442 924 646 1124
rect 498 706 590 924
rect 442 506 646 706
rect 498 474 590 506
rect 299 428 590 474
rect 500 366 510 369
rect 498 317 510 366
rect 578 366 588 369
rect 578 317 590 366
rect 498 288 590 317
rect 442 88 646 288
rect 301 7 311 59
rect 401 7 411 59
rect 498 10 590 88
rect 218 -31 276 -25
rect 218 -65 230 -31
rect 264 -65 276 -31
rect 218 -71 276 -65
<< via1 >>
rect 93 1571 183 1623
rect -84 1153 -16 1205
rect -84 425 -16 477
rect 93 7 183 59
rect 311 1571 401 1623
rect 510 1261 578 1313
rect 510 317 578 369
rect 311 7 401 59
<< metal2 >>
rect 93 1623 401 1633
rect 183 1571 311 1623
rect 93 1561 401 1571
rect 211 1313 578 1323
rect 211 1261 510 1313
rect 211 1251 578 1261
rect 211 1215 283 1251
rect -84 1205 283 1215
rect -16 1153 283 1205
rect -84 1143 283 1153
rect -84 477 283 487
rect -16 425 283 477
rect -84 415 283 425
rect 211 379 283 415
rect 211 369 578 379
rect 211 317 510 369
rect 211 307 578 317
rect 93 59 401 69
rect 183 7 311 59
rect 93 -3 401 7
use sky130_fd_pr__nfet_01v8_FZ7FED  sky130_fd_pr__nfet_01v8_FZ7FED_0
timestamp 1729325631
transform 1 0 247 0 1 815
box -247 -815 247 815
use sky130_fd_pr__nfet_01v8_V6EN4H  sky130_fd_pr__nfet_01v8_V6EN4H_0
timestamp 1729325631
transform 1 0 -50 0 1 815
box -108 -815 108 815
use sky130_fd_pr__nfet_01v8_V6EN4H  sky130_fd_pr__nfet_01v8_V6EN4H_1
timestamp 1729325631
transform 1 0 544 0 1 815
box -108 -815 108 815
<< labels >>
flabel poly 134 1434 134 1434 0 FreeSans 160 0 0 0 D6
port 0 nsew
flabel metal1 544 1454 544 1454 0 FreeSans 160 0 0 0 OUT
port 1 nsew
flabel metal1 246 1444 246 1444 0 FreeSans 160 0 0 0 GND
port 3 nsew
<< end >>
