magic
tech sky130A
magscale 1 2
timestamp 1729184099
<< error_p >>
rect -323 654 323 872
rect -323 18 323 236
rect -323 -618 323 -400
<< nwell >>
rect -323 654 323 1254
rect -323 18 323 618
rect -323 -618 323 -18
rect -323 -1254 323 -654
<< pmos >>
rect -229 754 -29 1154
rect 29 754 229 1154
rect -229 118 -29 518
rect 29 118 229 518
rect -229 -518 -29 -118
rect 29 -518 229 -118
rect -229 -1154 -29 -754
rect 29 -1154 229 -754
<< pdiff >>
rect -287 1142 -229 1154
rect -287 766 -275 1142
rect -241 766 -229 1142
rect -287 754 -229 766
rect -29 1142 29 1154
rect -29 766 -17 1142
rect 17 766 29 1142
rect -29 754 29 766
rect 229 1142 287 1154
rect 229 766 241 1142
rect 275 766 287 1142
rect 229 754 287 766
rect -287 506 -229 518
rect -287 130 -275 506
rect -241 130 -229 506
rect -287 118 -229 130
rect -29 506 29 518
rect -29 130 -17 506
rect 17 130 29 506
rect -29 118 29 130
rect 229 506 287 518
rect 229 130 241 506
rect 275 130 287 506
rect 229 118 287 130
rect -287 -130 -229 -118
rect -287 -506 -275 -130
rect -241 -506 -229 -130
rect -287 -518 -229 -506
rect -29 -130 29 -118
rect -29 -506 -17 -130
rect 17 -506 29 -130
rect -29 -518 29 -506
rect 229 -130 287 -118
rect 229 -506 241 -130
rect 275 -506 287 -130
rect 229 -518 287 -506
rect -287 -766 -229 -754
rect -287 -1142 -275 -766
rect -241 -1142 -229 -766
rect -287 -1154 -229 -1142
rect -29 -766 29 -754
rect -29 -1142 -17 -766
rect 17 -1142 29 -766
rect -29 -1154 29 -1142
rect 229 -766 287 -754
rect 229 -1142 241 -766
rect 275 -1142 287 -766
rect 229 -1154 287 -1142
<< pdiffc >>
rect -275 766 -241 1142
rect -17 766 17 1142
rect 241 766 275 1142
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
rect -275 -1142 -241 -766
rect -17 -1142 17 -766
rect 241 -1142 275 -766
<< poly >>
rect -229 1235 -29 1251
rect -229 1201 -213 1235
rect -45 1201 -29 1235
rect -229 1154 -29 1201
rect 29 1235 229 1251
rect 29 1201 45 1235
rect 213 1201 229 1235
rect 29 1154 229 1201
rect -229 707 -29 754
rect -229 673 -213 707
rect -45 673 -29 707
rect -229 657 -29 673
rect 29 707 229 754
rect 29 673 45 707
rect 213 673 229 707
rect 29 657 229 673
rect -229 599 -29 615
rect -229 565 -213 599
rect -45 565 -29 599
rect -229 518 -29 565
rect 29 599 229 615
rect 29 565 45 599
rect 213 565 229 599
rect 29 518 229 565
rect -229 71 -29 118
rect -229 37 -213 71
rect -45 37 -29 71
rect -229 21 -29 37
rect 29 71 229 118
rect 29 37 45 71
rect 213 37 229 71
rect 29 21 229 37
rect -229 -37 -29 -21
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect -229 -118 -29 -71
rect 29 -37 229 -21
rect 29 -71 45 -37
rect 213 -71 229 -37
rect 29 -118 229 -71
rect -229 -565 -29 -518
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect -229 -615 -29 -599
rect 29 -565 229 -518
rect 29 -599 45 -565
rect 213 -599 229 -565
rect 29 -615 229 -599
rect -229 -673 -29 -657
rect -229 -707 -213 -673
rect -45 -707 -29 -673
rect -229 -754 -29 -707
rect 29 -673 229 -657
rect 29 -707 45 -673
rect 213 -707 229 -673
rect 29 -754 229 -707
rect -229 -1201 -29 -1154
rect -229 -1235 -213 -1201
rect -45 -1235 -29 -1201
rect -229 -1251 -29 -1235
rect 29 -1201 229 -1154
rect 29 -1235 45 -1201
rect 213 -1235 229 -1201
rect 29 -1251 229 -1235
<< polycont >>
rect -213 1201 -45 1235
rect 45 1201 213 1235
rect -213 673 -45 707
rect 45 673 213 707
rect -213 565 -45 599
rect 45 565 213 599
rect -213 37 -45 71
rect 45 37 213 71
rect -213 -71 -45 -37
rect 45 -71 213 -37
rect -213 -599 -45 -565
rect 45 -599 213 -565
rect -213 -707 -45 -673
rect 45 -707 213 -673
rect -213 -1235 -45 -1201
rect 45 -1235 213 -1201
<< locali >>
rect -229 1201 -213 1235
rect -45 1201 -29 1235
rect 29 1201 45 1235
rect 213 1201 229 1235
rect -275 1142 -241 1158
rect -275 750 -241 766
rect -17 1142 17 1158
rect -17 750 17 766
rect 241 1142 275 1158
rect 241 750 275 766
rect -229 673 -213 707
rect -45 673 -29 707
rect 29 673 45 707
rect 213 673 229 707
rect -229 565 -213 599
rect -45 565 -29 599
rect 29 565 45 599
rect 213 565 229 599
rect -275 506 -241 522
rect -275 114 -241 130
rect -17 506 17 522
rect -17 114 17 130
rect 241 506 275 522
rect 241 114 275 130
rect -229 37 -213 71
rect -45 37 -29 71
rect 29 37 45 71
rect 213 37 229 71
rect -229 -71 -213 -37
rect -45 -71 -29 -37
rect 29 -71 45 -37
rect 213 -71 229 -37
rect -275 -130 -241 -114
rect -275 -522 -241 -506
rect -17 -130 17 -114
rect -17 -522 17 -506
rect 241 -130 275 -114
rect 241 -522 275 -506
rect -229 -599 -213 -565
rect -45 -599 -29 -565
rect 29 -599 45 -565
rect 213 -599 229 -565
rect -229 -707 -213 -673
rect -45 -707 -29 -673
rect 29 -707 45 -673
rect 213 -707 229 -673
rect -275 -766 -241 -750
rect -275 -1158 -241 -1142
rect -17 -766 17 -750
rect -17 -1158 17 -1142
rect 241 -766 275 -750
rect 241 -1158 275 -1142
rect -229 -1235 -213 -1201
rect -45 -1235 -29 -1201
rect 29 -1235 45 -1201
rect 213 -1235 229 -1201
<< viali >>
rect -192 1201 -66 1235
rect 66 1201 192 1235
rect -275 766 -241 1142
rect -17 766 17 1142
rect 241 766 275 1142
rect -192 673 -66 707
rect 66 673 192 707
rect -192 565 -66 599
rect 66 565 192 599
rect -275 130 -241 506
rect -17 130 17 506
rect 241 130 275 506
rect -192 37 -66 71
rect 66 37 192 71
rect -192 -71 -66 -37
rect 66 -71 192 -37
rect -275 -506 -241 -130
rect -17 -506 17 -130
rect 241 -506 275 -130
rect -192 -599 -66 -565
rect 66 -599 192 -565
rect -192 -707 -66 -673
rect 66 -707 192 -673
rect -275 -1142 -241 -766
rect -17 -1142 17 -766
rect 241 -1142 275 -766
rect -192 -1235 -66 -1201
rect 66 -1235 192 -1201
<< metal1 >>
rect -204 1235 -54 1241
rect -204 1201 -192 1235
rect -66 1201 -54 1235
rect -204 1195 -54 1201
rect 54 1235 204 1241
rect 54 1201 66 1235
rect 192 1201 204 1235
rect 54 1195 204 1201
rect -281 1142 -235 1154
rect -281 766 -275 1142
rect -241 766 -235 1142
rect -281 754 -235 766
rect -23 1142 23 1154
rect -23 766 -17 1142
rect 17 766 23 1142
rect -23 754 23 766
rect 235 1142 281 1154
rect 235 766 241 1142
rect 275 766 281 1142
rect 235 754 281 766
rect -204 707 -54 713
rect -204 673 -192 707
rect -66 673 -54 707
rect -204 667 -54 673
rect 54 707 204 713
rect 54 673 66 707
rect 192 673 204 707
rect 54 667 204 673
rect -204 599 -54 605
rect -204 565 -192 599
rect -66 565 -54 599
rect -204 559 -54 565
rect 54 599 204 605
rect 54 565 66 599
rect 192 565 204 599
rect 54 559 204 565
rect -281 506 -235 518
rect -281 130 -275 506
rect -241 130 -235 506
rect -281 118 -235 130
rect -23 506 23 518
rect -23 130 -17 506
rect 17 130 23 506
rect -23 118 23 130
rect 235 506 281 518
rect 235 130 241 506
rect 275 130 281 506
rect 235 118 281 130
rect -204 71 -54 77
rect -204 37 -192 71
rect -66 37 -54 71
rect -204 31 -54 37
rect 54 71 204 77
rect 54 37 66 71
rect 192 37 204 71
rect 54 31 204 37
rect -204 -37 -54 -31
rect -204 -71 -192 -37
rect -66 -71 -54 -37
rect -204 -77 -54 -71
rect 54 -37 204 -31
rect 54 -71 66 -37
rect 192 -71 204 -37
rect 54 -77 204 -71
rect -281 -130 -235 -118
rect -281 -506 -275 -130
rect -241 -506 -235 -130
rect -281 -518 -235 -506
rect -23 -130 23 -118
rect -23 -506 -17 -130
rect 17 -506 23 -130
rect -23 -518 23 -506
rect 235 -130 281 -118
rect 235 -506 241 -130
rect 275 -506 281 -130
rect 235 -518 281 -506
rect -204 -565 -54 -559
rect -204 -599 -192 -565
rect -66 -599 -54 -565
rect -204 -605 -54 -599
rect 54 -565 204 -559
rect 54 -599 66 -565
rect 192 -599 204 -565
rect 54 -605 204 -599
rect -204 -673 -54 -667
rect -204 -707 -192 -673
rect -66 -707 -54 -673
rect -204 -713 -54 -707
rect 54 -673 204 -667
rect 54 -707 66 -673
rect 192 -707 204 -673
rect 54 -713 204 -707
rect -281 -766 -235 -754
rect -281 -1142 -275 -766
rect -241 -1142 -235 -766
rect -281 -1154 -235 -1142
rect -23 -766 23 -754
rect -23 -1142 -17 -766
rect 17 -1142 23 -766
rect -23 -1154 23 -1142
rect 235 -766 281 -754
rect 235 -1142 241 -766
rect 275 -1142 281 -766
rect 235 -1154 281 -1142
rect -204 -1201 -54 -1195
rect -204 -1235 -192 -1201
rect -66 -1235 -54 -1201
rect -204 -1241 -54 -1235
rect 54 -1201 204 -1195
rect 54 -1235 66 -1201
rect 192 -1235 204 -1201
rect 54 -1241 204 -1235
<< properties >>
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 2 l 1 m 4 nf 2 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 75 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
