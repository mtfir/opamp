magic
tech sky130A
magscale 1 2
timestamp 1729217985
<< nmos >>
rect -41 109 41 509
rect -41 -509 41 -109
<< ndiff >>
rect -99 497 -41 509
rect -99 121 -87 497
rect -53 121 -41 497
rect -99 109 -41 121
rect 41 497 99 509
rect 41 121 53 497
rect 87 121 99 497
rect 41 109 99 121
rect -99 -121 -41 -109
rect -99 -497 -87 -121
rect -53 -497 -41 -121
rect -99 -509 -41 -497
rect 41 -121 99 -109
rect 41 -497 53 -121
rect 87 -497 99 -121
rect 41 -509 99 -497
<< ndiffc >>
rect -87 121 -53 497
rect 53 121 87 497
rect -87 -497 -53 -121
rect 53 -497 87 -121
<< poly >>
rect -41 581 41 597
rect -41 547 -25 581
rect 25 547 41 581
rect -41 509 41 547
rect -41 71 41 109
rect -41 37 -25 71
rect 25 37 41 71
rect -41 21 41 37
rect -41 -37 41 -21
rect -41 -71 -25 -37
rect 25 -71 41 -37
rect -41 -109 41 -71
rect -41 -547 41 -509
rect -41 -581 -25 -547
rect 25 -581 41 -547
rect -41 -597 41 -581
<< polycont >>
rect -25 547 25 581
rect -25 37 25 71
rect -25 -71 25 -37
rect -25 -581 25 -547
<< locali >>
rect -41 547 -25 581
rect 25 547 41 581
rect -87 497 -53 513
rect -87 105 -53 121
rect 53 497 87 513
rect 53 105 87 121
rect -41 37 -25 71
rect 25 37 41 71
rect -41 -71 -25 -37
rect 25 -71 41 -37
rect -87 -121 -53 -105
rect -87 -513 -53 -497
rect 53 -121 87 -105
rect 53 -513 87 -497
rect -41 -581 -25 -547
rect 25 -581 41 -547
<< viali >>
rect -25 547 25 581
rect -87 121 -53 497
rect 53 121 87 497
rect -25 37 25 71
rect -25 -71 25 -37
rect -87 -497 -53 -121
rect 53 -497 87 -121
rect -25 -581 25 -547
<< metal1 >>
rect -37 581 37 587
rect -37 547 -25 581
rect 25 547 37 581
rect -37 541 37 547
rect -93 497 -47 509
rect -93 121 -87 497
rect -53 121 -47 497
rect -93 109 -47 121
rect 47 497 93 509
rect 47 121 53 497
rect 87 121 93 497
rect 47 109 93 121
rect -37 71 37 77
rect -37 37 -25 71
rect 25 37 37 71
rect -37 31 37 37
rect -37 -37 37 -31
rect -37 -71 -25 -37
rect 25 -71 37 -37
rect -37 -77 37 -71
rect -93 -121 -47 -109
rect -93 -497 -87 -121
rect -53 -497 -47 -121
rect -93 -509 -47 -497
rect 47 -121 93 -109
rect 47 -497 53 -121
rect 87 -497 93 -121
rect 47 -509 93 -497
rect -37 -547 37 -541
rect -37 -581 -25 -547
rect 25 -581 37 -547
rect -37 -587 37 -581
<< properties >>
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 2 l 0.41 m 2 nf 1 diffcov 100 polycov 100 guard 0 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
