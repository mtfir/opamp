magic
tech sky130A
magscale 1 2
timestamp 1729411005
<< poly >>
rect 415 505 515 1335
rect 687 505 787 1335
<< viali >>
rect 573 1823 629 1857
rect 573 -17 629 17
<< metal1 >>
rect 561 1857 641 1863
rect 561 1823 573 1857
rect 629 1823 641 1857
rect 561 1817 641 1823
rect 147 1674 239 1761
rect 963 1674 1055 1761
rect 91 1474 409 1674
rect 521 1474 681 1674
rect 793 1474 1111 1674
rect 147 1436 239 1474
rect 147 1387 159 1436
rect 149 1384 159 1387
rect 227 1387 239 1436
rect 421 1433 431 1436
rect 419 1387 431 1433
rect 227 1384 237 1387
rect 421 1384 431 1387
rect 499 1433 509 1436
rect 499 1387 511 1433
rect 499 1384 509 1387
rect 149 1325 159 1328
rect 147 1276 159 1325
rect 227 1325 237 1328
rect 421 1325 431 1328
rect 227 1276 239 1325
rect 419 1279 431 1325
rect 421 1276 431 1279
rect 499 1325 509 1328
rect 499 1279 511 1325
rect 499 1276 509 1279
rect 147 1238 239 1276
rect 573 1238 629 1474
rect 963 1436 1055 1474
rect 693 1433 703 1436
rect 691 1387 703 1433
rect 693 1384 703 1387
rect 771 1433 781 1436
rect 771 1387 783 1433
rect 963 1387 975 1436
rect 771 1384 781 1387
rect 965 1384 975 1387
rect 1043 1387 1055 1436
rect 1043 1384 1053 1387
rect 693 1325 703 1328
rect 691 1279 703 1325
rect 693 1276 703 1279
rect 771 1325 781 1328
rect 965 1325 975 1328
rect 771 1279 783 1325
rect 771 1276 781 1279
rect 963 1276 975 1325
rect 1043 1325 1053 1328
rect 1043 1276 1055 1325
rect 963 1238 1055 1276
rect 91 1038 409 1238
rect 567 1038 635 1238
rect 793 1038 1111 1238
rect 147 802 239 1038
rect 573 802 629 1038
rect 963 802 1055 1038
rect 91 602 409 802
rect 567 602 635 802
rect 793 602 1111 802
rect 147 564 239 602
rect 147 515 159 564
rect 149 512 159 515
rect 227 515 239 564
rect 227 512 237 515
rect 421 512 431 564
rect 499 512 509 564
rect 149 453 159 456
rect 147 404 159 453
rect 227 453 237 456
rect 227 404 239 453
rect 421 404 431 456
rect 499 404 509 456
rect 147 366 239 404
rect 573 366 629 602
rect 963 564 1055 602
rect 693 512 703 564
rect 771 512 781 564
rect 963 515 975 564
rect 965 512 975 515
rect 1043 515 1055 564
rect 1043 512 1053 515
rect 693 404 703 456
rect 771 404 781 456
rect 965 453 975 456
rect 963 404 975 453
rect 1043 453 1053 456
rect 1043 404 1055 453
rect 963 366 1055 404
rect 91 166 409 366
rect 567 166 635 366
rect 793 166 1111 366
rect 147 79 239 166
rect 963 79 1055 166
rect 561 17 641 23
rect 561 -17 573 17
rect 629 -17 641 17
rect 561 -23 641 -17
<< via1 >>
rect 159 1384 227 1436
rect 431 1384 499 1436
rect 159 1276 227 1328
rect 431 1276 499 1328
rect 703 1384 771 1436
rect 975 1384 1043 1436
rect 703 1276 771 1328
rect 975 1276 1043 1328
rect 159 512 227 564
rect 431 512 499 564
rect 159 404 227 456
rect 431 404 499 456
rect 703 512 771 564
rect 975 512 1043 564
rect 703 404 771 456
rect 975 404 1043 456
<< metal2 >>
rect 21 1699 1181 1771
rect 21 1446 93 1699
rect 21 1436 227 1446
rect 21 1384 159 1436
rect 21 1374 227 1384
rect 431 1436 637 1446
rect 499 1384 637 1436
rect 431 1374 637 1384
rect 137 1336 248 1346
rect 137 1260 248 1270
rect 409 1335 521 1345
rect 409 1259 521 1269
rect 565 1338 637 1374
rect 681 1443 793 1453
rect 681 1367 793 1377
rect 953 1443 1065 1453
rect 953 1367 1065 1377
rect 1109 1338 1181 1699
rect 565 1328 771 1338
rect 565 1276 703 1328
rect 565 1266 771 1276
rect 975 1328 1181 1338
rect 1043 1276 1181 1328
rect 975 1266 1181 1276
rect 21 564 227 574
rect 21 512 159 564
rect 21 502 227 512
rect 431 564 637 574
rect 499 512 637 564
rect 431 502 637 512
rect 21 141 93 502
rect 137 458 249 473
rect 236 397 249 458
rect 137 387 249 397
rect 409 463 521 473
rect 409 387 521 397
rect 565 466 637 502
rect 681 571 793 581
rect 681 495 793 505
rect 953 566 1065 581
rect 1052 505 1065 566
rect 953 495 1065 505
rect 565 456 771 466
rect 565 404 703 456
rect 565 394 771 404
rect 975 456 1180 466
rect 1043 404 1180 456
rect 975 394 1180 404
rect 1108 141 1180 394
rect 21 69 1180 141
<< via2 >>
rect 137 1328 248 1336
rect 137 1276 159 1328
rect 159 1276 227 1328
rect 227 1276 248 1328
rect 137 1270 248 1276
rect 409 1328 521 1335
rect 409 1276 431 1328
rect 431 1276 499 1328
rect 499 1276 521 1328
rect 409 1269 521 1276
rect 681 1436 793 1443
rect 681 1384 703 1436
rect 703 1384 771 1436
rect 771 1384 793 1436
rect 681 1377 793 1384
rect 953 1436 1065 1443
rect 953 1384 975 1436
rect 975 1384 1043 1436
rect 1043 1384 1065 1436
rect 953 1377 1065 1384
rect 137 456 236 458
rect 137 404 159 456
rect 159 404 227 456
rect 227 404 236 456
rect 137 397 236 404
rect 409 456 521 463
rect 409 404 431 456
rect 431 404 499 456
rect 499 404 521 456
rect 409 397 521 404
rect 681 564 793 571
rect 681 512 703 564
rect 703 512 771 564
rect 771 512 793 564
rect 681 505 793 512
rect 953 564 1052 566
rect 953 512 975 564
rect 975 512 1043 564
rect 1043 512 1052 564
rect 953 505 1052 512
<< metal3 >>
rect 21 1695 1181 1771
rect 21 1341 97 1695
rect 1105 1448 1181 1695
rect 563 1443 803 1448
rect 563 1377 681 1443
rect 793 1377 803 1443
rect 563 1372 803 1377
rect 943 1443 1181 1448
rect 943 1377 953 1443
rect 1065 1377 1181 1443
rect 943 1372 1181 1377
rect 21 1336 258 1341
rect 563 1340 639 1372
rect 21 1270 137 1336
rect 248 1270 258 1336
rect 21 1265 258 1270
rect 399 1335 639 1340
rect 399 1269 409 1335
rect 521 1269 639 1335
rect 399 1264 639 1269
rect 563 571 803 576
rect 563 505 681 571
rect 793 505 803 571
rect 563 500 803 505
rect 932 566 1180 571
rect 932 505 953 566
rect 1052 505 1180 566
rect 563 468 639 500
rect 932 495 1180 505
rect 399 463 639 468
rect 21 458 248 463
rect 21 397 137 458
rect 236 397 248 458
rect 21 387 248 397
rect 399 397 409 463
rect 521 397 639 463
rect 399 392 639 397
rect 21 145 97 387
rect 1104 145 1180 495
rect 21 69 1180 145
use sky130_fd_pr__pfet_01v8_BHMD29  sky130_fd_pr__pfet_01v8_BHMD29_0
timestamp 1729312135
transform 1 0 601 0 1 920
box -654 -973 654 973
<< labels >>
flabel metal1 602 1570 602 1570 0 FreeSans 160 0 0 0 D5
port 0 nsew
flabel via1 466 1410 466 1410 0 FreeSans 160 0 0 0 VIN
port 1 nsew
flabel via2 740 1410 740 1410 0 FreeSans 160 0 0 0 VIP
port 2 nsew
flabel metal1 188 1577 188 1577 0 FreeSans 160 0 0 0 D6
port 3 nsew
flabel metal1 1011 1579 1011 1579 0 FreeSans 160 0 0 0 OUT
port 4 nsew
flabel viali 601 1842 601 1842 0 FreeSans 160 0 0 0 VDD
port 5 nsew
<< end >>
